module en_decode2_4 (out, enable, sel);
		output logic    [3:0] out;
		input logic     [1:0] sel;
		input logic        enable;
		
		